entity boxcar_filter is
  port (
    rst: in std_logic;
    clk: in std_logic;

    in_dat: in std_logic;
    in_clk: in std_logic;

    out
  ) ;
end boxcar_filter ;

architecture arch of boxcar_filter is



begin



end architecture ; -- arch